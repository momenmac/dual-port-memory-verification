class write_read_a_test extends test;
    function new(string name);
        super.new(name);
    endfunction

    virtual function void run();
        // Implement the test logic for write_read_a
    endfunction
endclass

class write_read_b_test extends test;
    function new(string name);
        super.new(name);
    endfunction

    virtual function void run();
        // Implement the test logic for write_read_b
    endfunction
endclass


class write_read_b_test extends test;
    function new(string name);
        super.new(name);
    endfunction

    virtual function void run();
        // Implement the test logic for write_read_b
    endfunction
endclass
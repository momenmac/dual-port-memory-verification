module tb;
    // Testbench code goes here
endmodule : tb
// Top-level testbench file that includes all components
`include "defines.sv"
`include "interface.sv"
`include "project_pkg.sv"
`include "../tests/basic_test.sv"
`include "../tests/extended_tests.sv"
`include "tb.sv"

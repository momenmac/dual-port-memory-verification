package project_pkg;
    // Include all the testbench components
    `include "transaction.sv"
    `include "test_registry.sv"
    `include "driver.sv"
//     `include "coverage.sv"
    `include "monitor.sv"
    `include "scoreboard.sv"
    `include "generator.sv"
    `include "agent.sv"
    `include "enviroment.sv"
endpackage

class write_read_a_generator extends generator;
    function new();
        super.new();
    endfunction

    virtual task run();
        // Implement specific logic for write_read_a test
        super.run();
    endtask

endclass


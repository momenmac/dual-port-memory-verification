class enviroment

endclass : enviroment
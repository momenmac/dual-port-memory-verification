class scoreboard;
    // scoreboard class to verify the correctness of transactions
endclass : scoreboard